library verilog;
use verilog.vl_types.all;
entity Checker_vlg_vec_tst is
end Checker_vlg_vec_tst;

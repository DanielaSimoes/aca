library verilog;
use verilog.vl_types.all;
entity Checker_vlg_check_tst is
    port(
        error           : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Checker_vlg_check_tst;

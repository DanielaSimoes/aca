library verilog;
use verilog.vl_types.all;
entity CRC_vlg_vec_tst is
end CRC_vlg_vec_tst;

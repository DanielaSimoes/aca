library verilog;
use verilog.vl_types.all;
entity ShiftRegister_vlg_vec_tst is
end ShiftRegister_vlg_vec_tst;
